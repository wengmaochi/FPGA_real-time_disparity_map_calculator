
module fp_qsys (
	altpll_100k_clk,
	altpll_100m_clk,
	altpll_100m_1_clk,
	altpll_12_5m_clk,
	altpll_25m_clk,
	clk_clk,
	reset_reset_n);	

	output		altpll_100k_clk;
	output		altpll_100m_clk;
	output		altpll_100m_1_clk;
	output		altpll_12_5m_clk;
	output		altpll_25m_clk;
	input		clk_clk;
	input		reset_reset_n;
endmodule

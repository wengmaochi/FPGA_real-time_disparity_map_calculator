    Mac OS X            	   2   �      �                                      ATTR       �   �   G                  �   G  com.apple.quarantine q/0081;61e2727e;Microsoft\x20Edge;F4DFF151-8F0D-4DA6-8F81-5C5FD694C068 